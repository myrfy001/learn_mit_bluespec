// TwoCycle.bsv
//
// This is a two cycle implementation of the RISC-V processor.

