// TwoStage.bsv
//
// This is a two stage pipelined implementation of the RISC-V processor.

